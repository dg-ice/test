module gdc_2020 (
input su;
output du;
);

endmodule
